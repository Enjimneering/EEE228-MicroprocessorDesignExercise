

module VGA_Driver (
    input wire        clk,
    input wire        reset,
    output reg        hsync,
    output reg        vsync,
    output reg  [9:0] x_pix,
    output reg  [9:0] y_pix
);








endmodule
