`ifndef SEG7MACROS
`define SEG7MACROS

`define CHAR_A 7'b0001000
`define CHAR_B 7'b0000011
`define CHAR_C 7'b1000110
`define CHAR_D 7'b0100001
`define CHAR_E 7'b0000110  
`define CHAR_F 7'b0001110  
`define CHAR_L 7'b1110001
`define CHAR_O 7'b1000000
`define CHAR_S 7'b0010010
`define CHAR_H 7'b0001001
`define CHAR_I 7'b0001001
`define CHAR_R 7'b1111010
`define CHAR_N 7'b1001001
`define CHAR_Z 7'b0100100
`define CHAR_U 7'b1000001
`define CHAR_P 7'b0001100
`define CHAR_T 7'b1110000
`define CHAR_V 7'b1000001  
`define CHAR_X 7'b0110000
`define CHAR_Y 7'b0010001
`define CHAR_ZERO 7'b1000000  
`define CHAR_ONE 7'b1111001  
`define CHAR_TWO  7'b0100100  
`define CHAR_THREE 7'b0110000  
`define CHAR_FOUR  7'b0011001  
`define CHAR_FIVE  7'b0010010  
`define CHAR_SIX   7'b0000010  
`define CHAR_SEVEN 7'b1111000  
`define CHAR_EIGHT 7'b0000000  
`define CHAR_NINE  7'b0010000  
`define CHAR_SPACE 7'b0010000  
      
`endif